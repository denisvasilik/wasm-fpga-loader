library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

package WasmFpgaLoaderPackage is

end package;

package body WasmFpgaLoaderPackage is

end package body;
